// Comprehensive Verilog version 7 exercise 15
// Template for shift-and-add multiplier exercise

`timescale 1ns / 1ns

module mult(
    input clk, reset,
    input [7:0] a, b,
    output [15:0] f,
    output busy
  );

endmodule
